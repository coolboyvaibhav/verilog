module Ripple_Add ();
    
    
endmodule